module aluf

import os
import net


fn build(){
        return $tmpl('../../../../../../../flag')
}
pub fn demo() {
        println(build())
}